module top (
	input clk,
	output [`LEDS_NR-1:0] led
);

reg [25:0] ctr_q;
wire [25:0] ctr_d;

// Sequential code (flip-flop)
always @(posedge clk)
	ctr_q <= ctr_d;

// Combinational code (boolean logic)
assign ctr_d = ctr_q + 1'b1;
assign led[`LEDS_NR-1:2] = {(`LEDS_NR - 2){1'b1}};
assign led[0] = ctr_q[25:25];

ODDR oddr_0(
	.D0(1'b0),
	.D1(1'b1),
	.CLK(ctr_q[25:25]),
	.Q0(led[1]),
	.Q1(),
	.TX(1'b0)
);

endmodule
