`default_nettype none

module top(output wire led);
	assign led = 1'b0;
endmodule

