`default_nettype none

module top(input wire resetn, output wire led);
	assign led = 1'b1;
endmodule

